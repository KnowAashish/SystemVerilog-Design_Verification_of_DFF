interface intf();

	bit		clk;
	logic 	resetn;
	logic 	din;
	logic 	dout;
	
endinterface