package dff_pkg;

`include "dff_transaction.sv"
`include "dff_generator.sv"
`include "dff_driver.sv"
`include "dff_monitor.sv"
`include "dff_scoreboard.sv"
`include "dff_env.sv"

endpackage